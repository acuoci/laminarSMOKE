THERMO ALL
300.   1000.   3500. 
H2                      H   2               G    300.00   3500.00  750.00      1
 3.73110902e+00-8.86706214e-04 1.12286897e-06-3.74349782e-10 4.17963674e-14    2
-1.08851547e+03-5.35285855e+00 3.08866003e+00 2.53968841e-03-5.72992027e-06    3
 5.71701843e-09-1.98865970e-12-9.92148124e+02-2.43823459e+00                   4
H2O                     H   2O   1          G    300.00   3500.00 1590.00      1
 2.30940463e+00 3.65433887e-03-1.22983871e-06 2.11931683e-10-1.50333493e-14    2
-2.97294901e+04 8.92765177e+00 4.03530937e+00-6.87559833e-04 2.86629214e-06    3
-1.50552360e-09 2.55006790e-13-3.02783278e+04-1.99201641e-01                   4
O2                      O   2               G    300.00   3500.00  760.00      1
 2.81750648e+00 2.49838007e-03-1.52493521e-06 4.50547608e-10-4.87702792e-14    2
-9.31713392e+02 7.94729337e+00 3.46035080e+00-8.85011121e-04 5.15281056e-06    3
-5.40712413e-09 1.87809542e-12-1.02942573e+03 5.02236126e+00                   4
N2                      N   2               G    300.00   3500.00 1050.00      1
 2.71287897e+00 1.90359754e-03-8.54297556e-07 1.84170938e-10-1.54715988e-14    2
-8.40225273e+02 7.15926558e+00 3.85321336e+00-2.44053349e-03 5.35160392e-06    3
-3.75608397e-09 9.22684330e-13-1.07969550e+03 1.60217419e+00                   4
END
