! This thermodynamic database was obtained by fitting the thermodynamic properties
! extracted from the following file: POLIMI_TOT_NOx_1407.CKT
! The thermodynamic properties are fitted in order to preserve not only the 
! continuity of each function at the intermediate temperature, but also the  continuity
! of the derivatives, from the 1st to the 3rd order
! The intermediate temperatures are chosen in order to minimize the fitting error.
! Last update: 1/20/2017

THERMO ALL
270.   1000.   3500. 
CH4                     C   1H   4          G    300.00   3500.00 1070.00      1
-2.82321418e-01 1.42739336e-02-6.77628877e-06 1.55380951e-09-1.39473841e-13    2
-9.36383584e+03 2.03507025e+01 2.85765313e+00 2.53571099e-03 9.67916347e-06    3
-8.69880871e-09 2.25599771e-12-1.00357904e+04 4.98969391e+00                   4
O2                      O   2               G    300.00   3500.00  760.00      1
 2.81750647e+00 2.49838008e-03-1.52493522e-06 4.50547610e-10-4.87702795e-14    2
-9.31713391e+02 7.94729338e+00 3.46035081e+00-8.85011180e-04 5.15281069e-06    3
-5.40712424e-09 1.87809546e-12-1.02942573e+03 5.02236122e+00                   4
CO2                     C   1O   2          G    300.00   3500.00 1620.00      1
 5.07830985e+00 2.05366041e-03-5.94311264e-07 5.38675127e-11 1.66346859e-15    2
-4.92442103e+04-4.47815291e+00 2.44892797e+00 8.54596135e-03-6.60570102e-06    3
 2.52769046e-09-3.80099332e-13-4.83922906e+04 9.47557732e+00                   4
CO                      C   1O   1          G    300.00   3500.00 1000.00      1
 2.68595014e+00 2.12486373e-03-1.04548609e-06 2.45538865e-10-2.22550982e-14    2
-1.41423615e+04 7.96579427e+00 3.81890943e+00-2.40697344e-03 5.75226967e-06    3
-4.28629830e-09 1.11070419e-12-1.43689533e+04 2.49992059e+00                   4
H2O                     H   2O   1          G    300.00   3500.00 1590.00      1
 2.30940463e+00 3.65433887e-03-1.22983871e-06 2.11931684e-10-1.50333493e-14    2
-2.97294901e+04 8.92765177e+00 4.03530937e+00-6.87559834e-04 2.86629215e-06    3
-1.50552360e-09 2.55006790e-13-3.02783278e+04-1.99201641e-01                   4
H2                      H   2               G    300.00   3500.00  750.00      1
 3.73110903e+00-8.86706228e-04 1.12286898e-06-3.74349786e-10 4.17963679e-14    2
-1.08851547e+03-5.35285858e+00 3.08866001e+00 2.53968852e-03-5.72992051e-06    3
 5.71701866e-09-1.98865978e-12-9.92148122e+02-2.43823451e+00                   4
H                       H   1               G    300.00   3500.00 1800.00      1
 2.50000000e+00-3.95459854e-15 2.96893838e-18-9.33318862e-22 1.04354326e-25    2
 2.54716200e+04-4.60117600e-01 2.50000000e+00 1.70660813e-16-4.68777753e-19    3
 3.39909334e-22-7.24829229e-26 2.54716200e+04-4.60117600e-01                   4
O                       O   1               G    300.00   3500.00  950.00      1
 2.57318360e+00-8.95609973e-05 4.05096293e-08-8.39812642e-12 9.43621954e-16    2
 2.92191409e+04 4.74952023e+00 2.95200330e+00-1.68459131e-03 2.55897855e-06    3
-1.77574473e-09 4.66034835e-13 2.91471652e+04 2.94136507e+00                   4
OH                      H   1O   1          G    300.00   3500.00  880.00      1
 3.62538437e+00-5.02165284e-04 8.36958465e-07-2.95714532e-10 3.30350487e-14    2
 3.41380110e+03 1.55419439e+00 3.37995108e+00 6.13440537e-04-1.06464237e-06    3
 1.14489216e-09-3.76228216e-13 3.45699735e+03 2.70689353e+00                   4
HO2                     H   1O   2          G    300.00   3500.00 1540.00      1
 4.16318067e+00 1.99798265e-03-4.89192085e-07 7.71153169e-11-7.30772101e-15    2
 4.41348946e+01 2.95517985e+00 2.85241381e+00 5.40257188e-03-3.80535043e-06    3
 1.51268170e-09-2.40354212e-13 4.47851086e+02 9.84483831e+00                   4
CH2                     C   1H   2          G    300.00   3500.00  900.00      1
 3.24505871e+00 2.75395076e-03-7.68471345e-07 8.23040044e-11-1.89900259e-15    2
 4.54794580e+04 4.28187007e+00 3.99717917e+00-5.88806836e-04 4.80279131e-06    3
-4.04455722e-09 1.14445134e-12 4.53440763e+04 7.32567425e-01                   4
CH2S                    C   1H   2          G    300.00   3500.00  900.00      1
 2.57518274e+00 4.11179660e-03-1.68232436e-06 3.44404950e-10-2.93085970e-14    2
 5.01958500e+04 6.99914505e+00 4.62572655e+00-5.00173142e-03 1.35068890e-05    3
-1.09068642e-08 3.09604395e-12 4.98267521e+04-2.67749713e+00                   4
CH3                     C   1H   3          G    300.00   3500.00 1270.00      1
 2.57723974e+00 6.62601164e-03-2.54906392e-06 4.67320141e-10-3.34867663e-14    2
 1.65488693e+04 6.94195966e+00 3.53327401e+00 3.61488008e-03 1.00739068e-06    3
-1.39958516e-09 3.34014278e-13 1.63060366e+04 2.10113860e+00                   4
HCO                     C   1H   1O   1     G    300.00   3500.00  920.00      1
 2.44772077e+00 5.65570556e-03-3.01329556e-06 7.57702525e-10-7.26129632e-14    2
 4.31149160e+03 1.15871953e+01 3.74218864e+00 2.75843940e-05 6.16298894e-06    3
-5.89177900e-09 1.73431136e-12 4.07330951e+03 5.45007089e+00                   4
CH2O                    C   1H   2O   1     G    300.00   3500.00  930.00      1
 1.06639253e+00 1.06960337e-02-5.54447373e-06 1.36053696e-09-1.28442555e-13    2
-1.46324373e+04 1.74071779e+01 3.13463322e+00 1.80037481e-03 8.80336319e-06    3
-8.92465079e-09 2.63639286e-12-1.50171301e+04 7.57920579e+00                   4
CH3OO                   C   1H   3O   2     G    300.00   3500.00 1300.00      1
 3.46521970e+00 1.23938518e-02-5.59614682e-06 1.22616716e-09-1.06238815e-13    2
 6.86982281e+02 1.04298931e+01 4.30117244e+00 9.82168948e-03-2.62826727e-06    3
-2.95822350e-10 1.86451475e-13 4.69634569e+02 6.17758023e+00                   4
C2H4                    C   2H   4          G    300.00   3500.00 1800.00      1
 4.49333672e+00 1.00335105e-02-3.62601388e-06 5.97613541e-10-3.65481279e-14    2
 3.93220822e+03-3.35192021e+00 2.66161697e-01 1.94272328e-02-1.14541158e-05    3
 3.49691054e-09-4.39228267e-13 5.45399123e+03 1.95264329e+01                   4
C2H5                    C   2H   5          G    300.00   3500.00  700.00      1
-1.10489358e+00 2.43511913e-02-1.39613152e-05 3.89870297e-09-4.17285120e-13    2
 1.35030749e+04 3.00146907e+01 4.99501829e+00-1.05054480e-02 6.07314832e-05    3
-6.72372955e-08 2.49884286e-11 1.26490872e+04 2.76182769e+00                   4
HCCO                    C   2H   1O   1     G    300.00   3500.00 1800.00      1
 7.44900313e+00 1.01177830e-03 3.02918166e-07-2.13909391e-10 2.81815209e-14    2
 1.86458955e+04-1.30987733e+01 4.44514163e+00 7.68702607e-03-5.25978830e-06    3
 1.84635226e-09-2.57965931e-13 1.97272856e+04 3.15875175e+00                   4
CH2CO                   C   2H   2O   1     G    300.00   3500.00 1410.00      1
 6.03578795e+00 5.81722421e-03-1.93206512e-06 2.83140053e-10-1.50051611e-14    2
-8.58422380e+03-7.64505060e+00 2.49197065e+00 1.58706066e-02-1.26271528e-05    3
 5.33991909e-09-9.11597189e-13-7.58486732e+03 1.06694385e+01                   4
CH2CHO                  C   2H   3O   1     G    300.00   3500.00 1030.00      1
 3.66502520e+00 1.44768244e-02-7.23266377e-06 1.70580456e-09-1.56345856e-13    2
-3.68579206e+01 5.92341848e+00 2.15742064e-01 2.78720987e-02-2.67403448e-05    3
 1.43321353e-08-3.22098925e-12 6.73694407e+02 2.26661724e+01                   4
C2H3                    C   2H   3          G    300.00   3500.00  700.00      1
 7.05094232e-01 1.53761148e-02-8.91788177e-06 2.51340904e-09-2.70561650e-13    2
 3.36189510e+04 1.96531878e+01 2.74606707e+00 3.71341285e-03 1.60736223e-05    3
-2.12880234e-08 8.22994995e-12 3.33332148e+04 1.05346375e+01                   4
C2H2                    C   2H   2          G    300.00   3500.00  970.00      1
 4.61193612e+00 5.01498203e-03-1.65253693e-06 2.49922529e-10-1.30568633e-14    2
 2.56043843e+04-3.75517098e+00 1.83812159e+00 1.64533925e-02-1.93408005e-05    3
 1.24068047e-08-3.14627392e-12 2.61425043e+04 9.54239254e+00                   4
N2                      N   2               G    300.00   3500.00 1050.00      1
 2.71287897e+00 1.90359754e-03-8.54297558e-07 1.84170938e-10-1.54715989e-14    2
-8.40225273e+02 7.15926558e+00 3.85321337e+00-2.44053350e-03 5.35160392e-06    3
-3.75608397e-09 9.22684332e-13-1.07969550e+03 1.60217419e+00                   4
END
